module top_module( 
    input [99:0] in,
    output [98:0] out_both,
    output [99:1] out_any,
    output [99:0] out_different );

for (integer i = 0; i < 99; i = i+1) begin
    
end

endmodule
